//======================================================================
//
// avalance_entropy.v
// ------------------
// Fake avalanche entropy source. This module SHOULD ONLY be used
// during simulation of the Cryptech True Random Number Generator
// (trng). The module DOES NOT provide any real entropy.
//
//
// Author: Joachim Strombergson
// Copyright (c) 2014, Secworks Sweden AB
// All rights reserved.
//
// Redistribution and use in source and binary forms, with or
// without modification, are permitted provided that the following
// conditions are met:
//
// 1. Redistributions of source code must retain the above copyright
//    notice, this list of conditions and the following disclaimer.
//
// 2. Redistributions in binary form must reproduce the above copyright
//    notice, this list of conditions and the following disclaimer in
//    the documentation and/or other materials provided with the
//    distribution.
//
// THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS
// "AS IS" AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT
// LIMITED TO, THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS
// FOR A PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
// COPYRIGHT OWNER OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT, INDIRECT,
// INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES (INCLUDING,
// BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES;
// LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER
// CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
// STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
// ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
// ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
//
//======================================================================

module avalance_entropy(
                        input wire           clk,
                        input wire           reset_n,

                        input wire           noise,

                        input wire           cs,
                        input wire           we,
                        input wire  [7 : 0]  address,
                        input wire  [31 : 0] write_data,
                        output wire [31 : 0] read_data,
                        output wire          error,

                        input wire           test_mode,
                        output wire          security_error,

                        output wire          entropy_enabled,
                        output wire [31 : 0] entropy_data,
                        output wire          entropy_valid,
                        input wire           entropy_ack,

                        output wire [7 : 0]  debug,
                        input wire           debug_update
                       );


  //----------------------------------------------------------------
  // Concurrent connectivity for ports etc.
  //----------------------------------------------------------------
  assign read_data      = 32'h00000000;
  assign error          = 0;
  assign security_error = 0;

  assign entropy_enabled = 1;
  assign entropy_data    = 32'h11223344;
  assign entropy_valid   = 1;

  assign debug           = 8'aa;

endmodule // avalance_entropy

//======================================================================
// EOF avalance_entropy.v
//======================================================================
